// Test top level design
`timescale 100 ps/ 100 ps

module test_top;

initial begin

    #1 $display("End of test");
end

endmodule
