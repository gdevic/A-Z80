// Copyright (C) 1991-2011 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 11.0 Build 208 07/03/2011 Service Pack 1 SJ Full Version"
// CREATED		"Mon Aug 18 07:13:24 2014"

module bus_control(
	ctl_bus_ff_oe,
	ctl_bus_zero_oe,
	ctl_bus_db_oe,
	bus_db_oe,
	db
);


input wire	ctl_bus_ff_oe;
input wire	ctl_bus_zero_oe;
input wire	ctl_bus_db_oe;
output wire	bus_db_oe;
inout wire	[7:0] db;

wire	[7:0] SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_5;
wire	[0:7] SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_4;

assign	SYNTHESIZED_WIRE_2 = 1;



assign	db[7] = SYNTHESIZED_WIRE_5 ? SYNTHESIZED_WIRE_0[7] : 1'bz;
assign	db[6] = SYNTHESIZED_WIRE_5 ? SYNTHESIZED_WIRE_0[6] : 1'bz;
assign	db[5] = SYNTHESIZED_WIRE_5 ? SYNTHESIZED_WIRE_0[5] : 1'bz;
assign	db[4] = SYNTHESIZED_WIRE_5 ? SYNTHESIZED_WIRE_0[4] : 1'bz;
assign	db[3] = SYNTHESIZED_WIRE_5 ? SYNTHESIZED_WIRE_0[3] : 1'bz;
assign	db[2] = SYNTHESIZED_WIRE_5 ? SYNTHESIZED_WIRE_0[2] : 1'bz;
assign	db[1] = SYNTHESIZED_WIRE_5 ? SYNTHESIZED_WIRE_0[1] : 1'bz;
assign	db[0] = SYNTHESIZED_WIRE_5 ? SYNTHESIZED_WIRE_0[0] : 1'bz;


assign	SYNTHESIZED_WIRE_0 = {ctl_bus_ff_oe,ctl_bus_ff_oe,ctl_bus_ff_oe,ctl_bus_ff_oe,ctl_bus_ff_oe,ctl_bus_ff_oe,ctl_bus_ff_oe,ctl_bus_ff_oe} & SYNTHESIZED_WIRE_2;

assign	SYNTHESIZED_WIRE_4 =  ~SYNTHESIZED_WIRE_5;

assign	bus_db_oe = ctl_bus_db_oe & SYNTHESIZED_WIRE_4;

assign	SYNTHESIZED_WIRE_5 = ctl_bus_ff_oe | ctl_bus_zero_oe;


endmodule
