// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
// CREATED		"Thu Dec 08 21:08:44 2016"

module resets(
	reset_in,
	clk,
	M1,
	T2,
	fpga_reset,
	hold_clk_wait,
	clrpc,
	nreset
);


input wire	reset_in;
input wire	clk;
input wire	M1;
input wire	T2;
input wire	fpga_reset;
input wire	hold_clk_wait;
output wire	clrpc;
output wire	nreset;

reg	clrpc_int;
wire	nclk;
reg	x1;
wire	x2;
wire	x3;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_1;
reg	SYNTHESIZED_WIRE_12;
reg	DFFE_intr_ff3;
reg	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_3;
reg	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_9;

assign	nreset = SYNTHESIZED_WIRE_9;




always@(posedge nclk or negedge SYNTHESIZED_WIRE_11)
begin
if (!SYNTHESIZED_WIRE_11)
	begin
	x1 <= 1;
	end
else
	begin
	x1 <= ~x1 & reset_in | x1 & ~SYNTHESIZED_WIRE_1;
	end
end

assign	clrpc = clrpc_int | SYNTHESIZED_WIRE_12 | DFFE_intr_ff3 | SYNTHESIZED_WIRE_13;

assign	SYNTHESIZED_WIRE_1 =  ~reset_in;

assign	x2 = x1 & SYNTHESIZED_WIRE_14;

assign	SYNTHESIZED_WIRE_14 = M1 & T2;

assign	x3 = x1 & SYNTHESIZED_WIRE_3;

assign	SYNTHESIZED_WIRE_9 =  ~SYNTHESIZED_WIRE_15;

assign	SYNTHESIZED_WIRE_16 =  ~hold_clk_wait;

assign	SYNTHESIZED_WIRE_3 =  ~SYNTHESIZED_WIRE_14;

assign	nclk =  ~clk;

assign	SYNTHESIZED_WIRE_11 =  ~fpga_reset;


always@(posedge nclk)
begin
if (SYNTHESIZED_WIRE_16)
	begin
	DFFE_intr_ff3 <= SYNTHESIZED_WIRE_12;
	end
end


always@(posedge nclk)
begin
if (SYNTHESIZED_WIRE_16)
	begin
	SYNTHESIZED_WIRE_13 <= SYNTHESIZED_WIRE_15;
	end
end


always@(posedge nclk)
begin
if (SYNTHESIZED_WIRE_16)
	begin
	SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_13;
	end
end


always@(posedge clk or negedge SYNTHESIZED_WIRE_11)
begin
if (!SYNTHESIZED_WIRE_11)
	begin
	SYNTHESIZED_WIRE_15 <= 1;
	end
else
	begin
	SYNTHESIZED_WIRE_15 <= x3;
	end
end


always@(posedge nclk or negedge SYNTHESIZED_WIRE_9)
begin
if (!SYNTHESIZED_WIRE_9)
	begin
	clrpc_int <= 0;
	end
else
	begin
	clrpc_int <= ~clrpc_int & x2 | clrpc_int & ~SYNTHESIZED_WIRE_14;
	end
end


endmodule
