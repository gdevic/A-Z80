//============================================================================
// Module execute in control/decode Z80 CPU
//
// Copyright 2014 Goran Devic
//
// This module implements the instruction execute state logic.
//============================================================================
`timescale 1ns/ 100 ps

module execute
(
    //----------------------------------------------------------
    // Control signals generated by the instruction execution
    //----------------------------------------------------------
    `include "exec_module.i"

    output logic nextM,
    output logic setM1,
    
    output logic fFetch,
    output logic fMRead,
    output logic fMWrite,
    output logic fIORead,
    output logic fIOWrite,
    
    output logic setM1ss,
    output logic setM1cc,
    output logic setM1bz,
    
    //----------------------------------------------------------
    // Inputs from the instruction decode PLA
    //----------------------------------------------------------
    input wire [104:0] pla,             // Statically decoded instructions

    //----------------------------------------------------------
    // Inputs from various blocks
    //----------------------------------------------------------
    input wire in_intr,                 // Servicing maskable interrupt
    input wire in_nmi,                  // Servicing non-maskable interrupt
    input wire im1,                     // Interrupt Mode 1
    input wire im2,                     // Interrupt Mode 2
    
    //----------------------------------------------------------
    // Machine and clock cycles
    //----------------------------------------------------------
    input wire M1,                      // Machine cycle #1
    input wire M2,                      // Machine cycle #2
    input wire M3,                      // Machine cycle #3
    input wire M4,                      // Machine cycle #4
    input wire M5,                      // Machine cycle #5
    input wire M6,                      // Machine cycle #6
    input wire T1,                      // T-cycle #1
    input wire T2,                      // T-cycle #2
    input wire T3,                      // T-cycle #3
    input wire T4,                      // T-cycle #4
    input wire T5,                      // T-cycle #5
    input wire T6                       // T-cycle #6
);

// If set by the execution matrix, prevents looping back to the next instruction
// Instructions that are longer than 4T set this at M1/T4
logic contM1;                           // Continue M1 cycle
// Instructions that use M2 immediately after M1/T4 set this at M1/T4
logic contM2;                           // Continue with the next M cycle

always_comb
begin
    contM1 = 0;
    contM2 = 0;

    //----------------------------------------------------------
    // Default assignment of all control outputs to 0 to prevent the
    // generation of latches
    //----------------------------------------------------------
    `include "exec_zero.i"

    //----------------------------------------------------------
    // State-based signal assignment
    //----------------------------------------------------------
    `include "exec_matrix.i"

    //----------------------------------------------------------
    // Default M1 fetch cycle execution
    //----------------------------------------------------------
    // M1 is a fetch phase
    if (M1) fFetch = 1;

    if (M1 && T1) begin     // T1: PC => AB
        ctl_reg_sel_pc = 1;
        ctl_al_we = 1;
    end
    
    if (M1 && T2) begin     // T2: Incr(PC); Get opcode from DB
    
        ctl_ir_we = 1;
        ctl_bus_inc_we = 1;
        
        // When servicing interrupts, depending on the interrupt mode:
        // IM0 : (nothing special here)
        // IM1 : Force FF on the bus and execute it (RST38 instruction)
        // IM2 : Force 00 on the bus - later we execute a special CALL on that NOP
        // NMI : Force FF on the bus and execute it (RST38 instruction)
        //       within the RST instruction the target address is conditionally set to 0x66
        if (in_intr || in_nmi) begin
            if (in_intr) begin
                if (im1) ctl_bus_ff_oe = 1;
                if (im2) ctl_bus_zero_oe = 1;
            end else    // in_nmi
                ctl_bus_ff_oe = 1;
        end else begin
            ctl_bus_db_oe = 1;
        end
    end

    if (M1 && T3) begin
    end

    // At T4, evaluate continuation flags for some instructions that need more than 4T
    if (M1 && T4) begin
        nextM = !contM1;
        setM1 = !contM1 & !contM2;
    end

end

endmodule
